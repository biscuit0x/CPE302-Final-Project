library verilog;
use verilog.vl_types.all;
entity TOP_vlg_sample_tst is
    port(
        CLK             : in     vl_logic;
        RESET           : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end TOP_vlg_sample_tst;
